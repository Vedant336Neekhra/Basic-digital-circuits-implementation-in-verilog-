module demo();

    initial
    begin
      $display("hello ,world");
    end

endmodule